module counter_scratch#(
    //parameter
    parameter WIDTH = 1
)(
    //input
    input wire rst,
    input wire clk,
    //output
    output wire [0:WIDTH-1] count
);
endmodule

